module subtractor(
  input in1,
  input in2,
  output out)

  out = in1 - in2

endmodule
